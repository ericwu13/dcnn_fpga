// qsysP01_tb.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module qsysP01_tb (
	);

	wire         qsysp01_inst_clk_bfm_clk_clk;          // qsysP01_inst_clk_bfm:clk -> [qsysP01_inst:clk_clk, qsysP01_inst_reset_bfm:clk]
	wire   [6:0] qsysp01_inst_hex_out_export;           // qsysP01_inst:hex_out_export -> qsysP01_inst_hex_out_bfm:sig_export
	wire  [17:0] qsysp01_inst_led_out_export;           // qsysP01_inst:led_out_export -> qsysP01_inst_led_out_bfm:sig_export
	wire         qsysp01_inst_rs232_ex_txd;             // qsysP01_inst:rs232_ex_TXD -> qsysP01_inst_rs232_ex_bfm:sig_TXD
	wire   [0:0] qsysp01_inst_rs232_ex_bfm_conduit_rxd; // qsysP01_inst_rs232_ex_bfm:sig_RXD -> qsysP01_inst:rs232_ex_RXD
	wire         qsysp01_inst_sdram_w_cs_n;             // qsysP01_inst:sdram_w_cs_n -> qsysP01_inst_sdram_w_bfm:sig_cs_n
	wire   [3:0] qsysp01_inst_sdram_w_dqm;              // qsysP01_inst:sdram_w_dqm -> qsysP01_inst_sdram_w_bfm:sig_dqm
	wire         qsysp01_inst_sdram_w_cas_n;            // qsysP01_inst:sdram_w_cas_n -> qsysP01_inst_sdram_w_bfm:sig_cas_n
	wire         qsysp01_inst_sdram_w_ras_n;            // qsysP01_inst:sdram_w_ras_n -> qsysP01_inst_sdram_w_bfm:sig_ras_n
	wire         qsysp01_inst_sdram_w_we_n;             // qsysP01_inst:sdram_w_we_n -> qsysP01_inst_sdram_w_bfm:sig_we_n
	wire  [12:0] qsysp01_inst_sdram_w_addr;             // qsysP01_inst:sdram_w_addr -> qsysP01_inst_sdram_w_bfm:sig_addr
	wire         qsysp01_inst_sdram_w_cke;              // qsysP01_inst:sdram_w_cke -> qsysP01_inst_sdram_w_bfm:sig_cke
	wire  [31:0] qsysp01_inst_sdram_w_dq;               // [] -> [qsysP01_inst:sdram_w_dq, qsysP01_inst_sdram_w_bfm:sig_dq]
	wire   [1:0] qsysp01_inst_sdram_w_ba;               // qsysP01_inst:sdram_w_ba -> qsysP01_inst_sdram_w_bfm:sig_ba
	wire  [17:0] qsysp01_inst_sw_in_bfm_conduit_export; // qsysP01_inst_sw_in_bfm:sig_export -> qsysP01_inst:sw_in_export
	wire         qsysp01_inst_reset_bfm_reset_reset;    // qsysP01_inst_reset_bfm:reset -> qsysP01_inst:reset_reset_n

	qsysP01 qsysp01_inst (
		.clk_clk        (qsysp01_inst_clk_bfm_clk_clk),          //       clk.clk
		.hex_out_export (qsysp01_inst_hex_out_export),           //   hex_out.export
		.led_out_export (qsysp01_inst_led_out_export),           //   led_out.export
		.reset_reset_n  (qsysp01_inst_reset_bfm_reset_reset),    //     reset.reset_n
		.rs232_ex_RXD   (qsysp01_inst_rs232_ex_bfm_conduit_rxd), //  rs232_ex.RXD
		.rs232_ex_TXD   (qsysp01_inst_rs232_ex_txd),             //          .TXD
		.sdram_clk_clk  (),                                      // sdram_clk.clk
		.sdram_w_addr   (qsysp01_inst_sdram_w_addr),             //   sdram_w.addr
		.sdram_w_ba     (qsysp01_inst_sdram_w_ba),               //          .ba
		.sdram_w_cas_n  (qsysp01_inst_sdram_w_cas_n),            //          .cas_n
		.sdram_w_cke    (qsysp01_inst_sdram_w_cke),              //          .cke
		.sdram_w_cs_n   (qsysp01_inst_sdram_w_cs_n),             //          .cs_n
		.sdram_w_dq     (qsysp01_inst_sdram_w_dq),               //          .dq
		.sdram_w_dqm    (qsysp01_inst_sdram_w_dqm),              //          .dqm
		.sdram_w_ras_n  (qsysp01_inst_sdram_w_ras_n),            //          .ras_n
		.sdram_w_we_n   (qsysp01_inst_sdram_w_we_n),             //          .we_n
		.sw_in_export   (qsysp01_inst_sw_in_bfm_conduit_export)  //     sw_in.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) qsysp01_inst_clk_bfm (
		.clk (qsysp01_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm qsysp01_inst_hex_out_bfm (
		.sig_export (qsysp01_inst_hex_out_export)  // conduit.export
	);

	altera_conduit_bfm_0002 qsysp01_inst_led_out_bfm (
		.sig_export (qsysp01_inst_led_out_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) qsysp01_inst_reset_bfm (
		.reset (qsysp01_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (qsysp01_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 qsysp01_inst_rs232_ex_bfm (
		.sig_RXD (qsysp01_inst_rs232_ex_bfm_conduit_rxd), // conduit.RXD
		.sig_TXD (qsysp01_inst_rs232_ex_txd)              //        .TXD
	);

	altera_conduit_bfm_0004 qsysp01_inst_sdram_w_bfm (
		.sig_addr  (qsysp01_inst_sdram_w_addr),  // conduit.addr
		.sig_ba    (qsysp01_inst_sdram_w_ba),    //        .ba
		.sig_cas_n (qsysp01_inst_sdram_w_cas_n), //        .cas_n
		.sig_cke   (qsysp01_inst_sdram_w_cke),   //        .cke
		.sig_cs_n  (qsysp01_inst_sdram_w_cs_n),  //        .cs_n
		.sig_dq    (qsysp01_inst_sdram_w_dq),    //        .dq
		.sig_dqm   (qsysp01_inst_sdram_w_dqm),   //        .dqm
		.sig_ras_n (qsysp01_inst_sdram_w_ras_n), //        .ras_n
		.sig_we_n  (qsysp01_inst_sdram_w_we_n)   //        .we_n
	);

	altera_conduit_bfm_0005 qsysp01_inst_sw_in_bfm (
		.sig_export (qsysp01_inst_sw_in_bfm_conduit_export)  // conduit.export
	);

endmodule
