// qsysP01.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module qsysP01 (
		input  wire        clk_clk,        //       clk.clk
		output wire [6:0]  hex_out_export, //   hex_out.export
		output wire [17:0] led_out_export, //   led_out.export
		input  wire        reset_reset_n,  //     reset.reset_n
		input  wire        rs232_ex_RXD,   //  rs232_ex.RXD
		output wire        rs232_ex_TXD,   //          .TXD
		output wire        sdram_clk_clk,  // sdram_clk.clk
		output wire [12:0] sdram_w_addr,   //   sdram_w.addr
		output wire [1:0]  sdram_w_ba,     //          .ba
		output wire        sdram_w_cas_n,  //          .cas_n
		output wire        sdram_w_cke,    //          .cke
		output wire        sdram_w_cs_n,   //          .cs_n
		inout  wire [31:0] sdram_w_dq,     //          .dq
		output wire [3:0]  sdram_w_dqm,    //          .dqm
		output wire        sdram_w_ras_n,  //          .ras_n
		output wire        sdram_w_we_n,   //          .we_n
		input  wire [17:0] sw_in_export    //     sw_in.export
	);

	wire         altpll_0_c1_clk;                                             // altpll_0:c1 -> [hex0_output:clk, irq_mapper:clk, jtag_uart_0:clk, led_output:clk, mm_interconnect_0:altpll_0_c1_clk, nios2:clk, onchip_memory2_0:clk, rs232_0:clk, rst_controller_001:clk, sdram_control:clk, sw_input:clk, sysid_qsys_0:clock, test_slave_0:i_clk_ctrl]
	wire  [31:0] nios2_data_master_readdata;                                  // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                               // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                               // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [28:0] nios2_data_master_address;                                   // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                      // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_readdatavalid;                             // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire         nios2_data_master_write;                                     // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                 // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                           // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [28:0] nios2_instruction_master_address;                            // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                               // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect;     // mm_interconnect_0:rs232_0_avalon_rs232_slave_chipselect -> rs232_0:chipselect
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata;       // rs232_0:readdata -> mm_interconnect_0:rs232_0_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_address;        // mm_interconnect_0:rs232_0_avalon_rs232_slave_address -> rs232_0:address
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_read;           // mm_interconnect_0:rs232_0_avalon_rs232_slave_read -> rs232_0:read
	wire   [3:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable;     // mm_interconnect_0:rs232_0_avalon_rs232_slave_byteenable -> rs232_0:byteenable
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_write;          // mm_interconnect_0:rs232_0_avalon_rs232_slave_write -> rs232_0:write
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata;      // mm_interconnect_0:rs232_0_avalon_rs232_slave_writedata -> rs232_0:writedata
	wire  [31:0] mm_interconnect_0_test_slave_0_avalon_slave_0_readdata;      // test_slave_0:o_y_data -> mm_interconnect_0:test_slave_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_test_slave_0_avalon_slave_0_waitrequest;   // test_slave_0:o_wait_req -> mm_interconnect_0:test_slave_0_avalon_slave_0_waitrequest
	wire         mm_interconnect_0_test_slave_0_avalon_slave_0_read;          // mm_interconnect_0:test_slave_0_avalon_slave_0_read -> test_slave_0:i_read_req
	wire         mm_interconnect_0_test_slave_0_avalon_slave_0_write;         // mm_interconnect_0:test_slave_0_avalon_slave_0_write -> test_slave_0:i_write_req
	wire  [31:0] mm_interconnect_0_test_slave_0_avalon_slave_0_writedata;     // mm_interconnect_0:test_slave_0_avalon_slave_0_writedata -> test_slave_0:i_data_32b_ctrl
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;            // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;         // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;             // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;               // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;               // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                   // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                  // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;              // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_sdram_control_s1_chipselect;               // mm_interconnect_0:sdram_control_s1_chipselect -> sdram_control:az_cs
	wire  [31:0] mm_interconnect_0_sdram_control_s1_readdata;                 // sdram_control:za_data -> mm_interconnect_0:sdram_control_s1_readdata
	wire         mm_interconnect_0_sdram_control_s1_waitrequest;              // sdram_control:za_waitrequest -> mm_interconnect_0:sdram_control_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_control_s1_address;                  // mm_interconnect_0:sdram_control_s1_address -> sdram_control:az_addr
	wire         mm_interconnect_0_sdram_control_s1_read;                     // mm_interconnect_0:sdram_control_s1_read -> sdram_control:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_control_s1_byteenable;               // mm_interconnect_0:sdram_control_s1_byteenable -> sdram_control:az_be_n
	wire         mm_interconnect_0_sdram_control_s1_readdatavalid;            // sdram_control:za_valid -> mm_interconnect_0:sdram_control_s1_readdatavalid
	wire         mm_interconnect_0_sdram_control_s1_write;                    // mm_interconnect_0:sdram_control_s1_write -> sdram_control:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_control_s1_writedata;                // mm_interconnect_0:sdram_control_s1_writedata -> sdram_control:az_data
	wire  [31:0] mm_interconnect_0_sw_input_s1_readdata;                      // sw_input:readdata -> mm_interconnect_0:sw_input_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_input_s1_address;                       // mm_interconnect_0:sw_input_s1_address -> sw_input:address
	wire         mm_interconnect_0_led_output_s1_chipselect;                  // mm_interconnect_0:led_output_s1_chipselect -> led_output:chipselect
	wire  [31:0] mm_interconnect_0_led_output_s1_readdata;                    // led_output:readdata -> mm_interconnect_0:led_output_s1_readdata
	wire   [1:0] mm_interconnect_0_led_output_s1_address;                     // mm_interconnect_0:led_output_s1_address -> led_output:address
	wire         mm_interconnect_0_led_output_s1_write;                       // mm_interconnect_0:led_output_s1_write -> led_output:write_n
	wire  [31:0] mm_interconnect_0_led_output_s1_writedata;                   // mm_interconnect_0:led_output_s1_writedata -> led_output:writedata
	wire         mm_interconnect_0_hex0_output_s1_chipselect;                 // mm_interconnect_0:hex0_output_s1_chipselect -> hex0_output:chipselect
	wire  [31:0] mm_interconnect_0_hex0_output_s1_readdata;                   // hex0_output:readdata -> mm_interconnect_0:hex0_output_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_output_s1_address;                    // mm_interconnect_0:hex0_output_s1_address -> hex0_output:address
	wire         mm_interconnect_0_hex0_output_s1_write;                      // mm_interconnect_0:hex0_output_s1_write -> hex0_output:write_n
	wire  [31:0] mm_interconnect_0_hex0_output_s1_writedata;                  // mm_interconnect_0:hex0_output_s1_writedata -> hex0_output:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [16:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // rs232_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                               // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         nios2_debug_reset_request_reset;                             // nios2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [hex0_output:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, led_output:reset_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, onchip_memory2_0:reset, rs232_0:reset, rst_translator:in_reset, sdram_control:reset_n, sw_input:reset_n, sysid_qsys_0:reset_n, test_slave_0:i_rst_ctrl]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	qsysP01_altpll_0 altpll_0 (
		.clk       (clk_clk),                                        //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0        (sdram_clk_clk),                                  //                    c0.clk
		.c1        (altpll_0_c1_clk),                                //                    c1.clk
		.areset    (),                                               //        areset_conduit.export
		.locked    (),                                               //        locked_conduit.export
		.phasedone ()                                                //     phasedone_conduit.export
	);

	qsysP01_hex0_output hex0_output (
		.clk        (altpll_0_c1_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_hex0_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_output_s1_readdata),   //                    .readdata
		.out_port   (hex_out_export)                               // external_connection.export
	);

	qsysP01_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c1_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	qsysP01_led_output led_output (
		.clk        (altpll_0_c1_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_led_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_output_s1_readdata),   //                    .readdata
		.out_port   (led_out_export)                              // external_connection.export
	);

	qsysP01_nios2 nios2 (
		.clk                                 (altpll_0_c1_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	qsysP01_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c1_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	qsysP01_rs232_0 rs232_0 (
		.clk        (altpll_0_c1_clk),                                         //                clk.clk
		.reset      (rst_controller_001_reset_out_reset),                      //              reset.reset
		.address    (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                                //          interrupt.irq
		.UART_RXD   (rs232_ex_RXD),                                            // external_interface.export
		.UART_TXD   (rs232_ex_TXD)                                             //                   .export
	);

	qsysP01_sdram_control sdram_control (
		.clk            (altpll_0_c1_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),              // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_control_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_control_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_control_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_control_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_control_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_control_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_control_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_control_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_control_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_w_addr),                                     //  wire.export
		.zs_ba          (sdram_w_ba),                                       //      .export
		.zs_cas_n       (sdram_w_cas_n),                                    //      .export
		.zs_cke         (sdram_w_cke),                                      //      .export
		.zs_cs_n        (sdram_w_cs_n),                                     //      .export
		.zs_dq          (sdram_w_dq),                                       //      .export
		.zs_dqm         (sdram_w_dqm),                                      //      .export
		.zs_ras_n       (sdram_w_ras_n),                                    //      .export
		.zs_we_n        (sdram_w_we_n)                                      //      .export
	);

	qsysP01_sw_input sw_input (
		.clk      (altpll_0_c1_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_sw_input_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_input_s1_readdata), //                    .readdata
		.in_port  (sw_in_export)                            // external_connection.export
	);

	qsysP01_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c1_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	qsysP01_test_slave_0 test_slave_0 (
		.i_data_32b_ctrl (mm_interconnect_0_test_slave_0_avalon_slave_0_writedata),   // avalon_slave_0.writedata
		.o_wait_req      (mm_interconnect_0_test_slave_0_avalon_slave_0_waitrequest), //               .waitrequest
		.o_y_data        (mm_interconnect_0_test_slave_0_avalon_slave_0_readdata),    //               .readdata
		.i_read_req      (mm_interconnect_0_test_slave_0_avalon_slave_0_read),        //               .read
		.i_write_req     (mm_interconnect_0_test_slave_0_avalon_slave_0_write),       //               .write
		.i_clk_ctrl      (altpll_0_c1_clk),                                           //     clock_sink.clk
		.i_rst_ctrl      (rst_controller_001_reset_out_reset)                         //     reset_sink.reset
	);

	qsysP01_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c1_clk                                            (altpll_0_c1_clk),                                             //                                          altpll_0_c1.clk
		.clk_0_clk_clk                                              (clk_clk),                                                     //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_reset_reset_bridge_in_reset_reset                    (rst_controller_001_reset_out_reset),                          //                    nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                                  (nios2_data_master_address),                                   //                                    nios2_data_master.address
		.nios2_data_master_waitrequest                              (nios2_data_master_waitrequest),                               //                                                     .waitrequest
		.nios2_data_master_byteenable                               (nios2_data_master_byteenable),                                //                                                     .byteenable
		.nios2_data_master_read                                     (nios2_data_master_read),                                      //                                                     .read
		.nios2_data_master_readdata                                 (nios2_data_master_readdata),                                  //                                                     .readdata
		.nios2_data_master_readdatavalid                            (nios2_data_master_readdatavalid),                             //                                                     .readdatavalid
		.nios2_data_master_write                                    (nios2_data_master_write),                                     //                                                     .write
		.nios2_data_master_writedata                                (nios2_data_master_writedata),                                 //                                                     .writedata
		.nios2_data_master_debugaccess                              (nios2_data_master_debugaccess),                               //                                                     .debugaccess
		.nios2_instruction_master_address                           (nios2_instruction_master_address),                            //                             nios2_instruction_master.address
		.nios2_instruction_master_waitrequest                       (nios2_instruction_master_waitrequest),                        //                                                     .waitrequest
		.nios2_instruction_master_read                              (nios2_instruction_master_read),                               //                                                     .read
		.nios2_instruction_master_readdata                          (nios2_instruction_master_readdata),                           //                                                     .readdata
		.nios2_instruction_master_readdatavalid                     (nios2_instruction_master_readdatavalid),                      //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                  //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                   //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),               //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),              //                                                     .writedata
		.hex0_output_s1_address                                     (mm_interconnect_0_hex0_output_s1_address),                    //                                       hex0_output_s1.address
		.hex0_output_s1_write                                       (mm_interconnect_0_hex0_output_s1_write),                      //                                                     .write
		.hex0_output_s1_readdata                                    (mm_interconnect_0_hex0_output_s1_readdata),                   //                                                     .readdata
		.hex0_output_s1_writedata                                   (mm_interconnect_0_hex0_output_s1_writedata),                  //                                                     .writedata
		.hex0_output_s1_chipselect                                  (mm_interconnect_0_hex0_output_s1_chipselect),                 //                                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                     .chipselect
		.led_output_s1_address                                      (mm_interconnect_0_led_output_s1_address),                     //                                        led_output_s1.address
		.led_output_s1_write                                        (mm_interconnect_0_led_output_s1_write),                       //                                                     .write
		.led_output_s1_readdata                                     (mm_interconnect_0_led_output_s1_readdata),                    //                                                     .readdata
		.led_output_s1_writedata                                    (mm_interconnect_0_led_output_s1_writedata),                   //                                                     .writedata
		.led_output_s1_chipselect                                   (mm_interconnect_0_led_output_s1_chipselect),                  //                                                     .chipselect
		.nios2_debug_mem_slave_address                              (mm_interconnect_0_nios2_debug_mem_slave_address),             //                                nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                                (mm_interconnect_0_nios2_debug_mem_slave_write),               //                                                     .write
		.nios2_debug_mem_slave_read                                 (mm_interconnect_0_nios2_debug_mem_slave_read),                //                                                     .read
		.nios2_debug_mem_slave_readdata                             (mm_interconnect_0_nios2_debug_mem_slave_readdata),            //                                                     .readdata
		.nios2_debug_mem_slave_writedata                            (mm_interconnect_0_nios2_debug_mem_slave_writedata),           //                                                     .writedata
		.nios2_debug_mem_slave_byteenable                           (mm_interconnect_0_nios2_debug_mem_slave_byteenable),          //                                                     .byteenable
		.nios2_debug_mem_slave_waitrequest                          (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),         //                                                     .waitrequest
		.nios2_debug_mem_slave_debugaccess                          (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),         //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),               //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                                     .clken
		.rs232_0_avalon_rs232_slave_address                         (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),        //                           rs232_0_avalon_rs232_slave.address
		.rs232_0_avalon_rs232_slave_write                           (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),          //                                                     .write
		.rs232_0_avalon_rs232_slave_read                            (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),           //                                                     .read
		.rs232_0_avalon_rs232_slave_readdata                        (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),       //                                                     .readdata
		.rs232_0_avalon_rs232_slave_writedata                       (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),      //                                                     .writedata
		.rs232_0_avalon_rs232_slave_byteenable                      (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable),     //                                                     .byteenable
		.rs232_0_avalon_rs232_slave_chipselect                      (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect),     //                                                     .chipselect
		.sdram_control_s1_address                                   (mm_interconnect_0_sdram_control_s1_address),                  //                                     sdram_control_s1.address
		.sdram_control_s1_write                                     (mm_interconnect_0_sdram_control_s1_write),                    //                                                     .write
		.sdram_control_s1_read                                      (mm_interconnect_0_sdram_control_s1_read),                     //                                                     .read
		.sdram_control_s1_readdata                                  (mm_interconnect_0_sdram_control_s1_readdata),                 //                                                     .readdata
		.sdram_control_s1_writedata                                 (mm_interconnect_0_sdram_control_s1_writedata),                //                                                     .writedata
		.sdram_control_s1_byteenable                                (mm_interconnect_0_sdram_control_s1_byteenable),               //                                                     .byteenable
		.sdram_control_s1_readdatavalid                             (mm_interconnect_0_sdram_control_s1_readdatavalid),            //                                                     .readdatavalid
		.sdram_control_s1_waitrequest                               (mm_interconnect_0_sdram_control_s1_waitrequest),              //                                                     .waitrequest
		.sdram_control_s1_chipselect                                (mm_interconnect_0_sdram_control_s1_chipselect),               //                                                     .chipselect
		.sw_input_s1_address                                        (mm_interconnect_0_sw_input_s1_address),                       //                                          sw_input_s1.address
		.sw_input_s1_readdata                                       (mm_interconnect_0_sw_input_s1_readdata),                      //                                                     .readdata
		.sysid_qsys_0_control_slave_address                         (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //                           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                                     .readdata
		.test_slave_0_avalon_slave_0_write                          (mm_interconnect_0_test_slave_0_avalon_slave_0_write),         //                          test_slave_0_avalon_slave_0.write
		.test_slave_0_avalon_slave_0_read                           (mm_interconnect_0_test_slave_0_avalon_slave_0_read),          //                                                     .read
		.test_slave_0_avalon_slave_0_readdata                       (mm_interconnect_0_test_slave_0_avalon_slave_0_readdata),      //                                                     .readdata
		.test_slave_0_avalon_slave_0_writedata                      (mm_interconnect_0_test_slave_0_avalon_slave_0_writedata),     //                                                     .writedata
		.test_slave_0_avalon_slave_0_waitrequest                    (mm_interconnect_0_test_slave_0_avalon_slave_0_waitrequest)    //                                                     .waitrequest
	);

	qsysP01_irq_mapper irq_mapper (
		.clk           (altpll_0_c1_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                  // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                // (terminated)
		.reset_req_in0  (1'b0),                            // (terminated)
		.reset_req_in1  (1'b0),                            // (terminated)
		.reset_in2      (1'b0),                            // (terminated)
		.reset_req_in2  (1'b0),                            // (terminated)
		.reset_in3      (1'b0),                            // (terminated)
		.reset_req_in3  (1'b0),                            // (terminated)
		.reset_in4      (1'b0),                            // (terminated)
		.reset_req_in4  (1'b0),                            // (terminated)
		.reset_in5      (1'b0),                            // (terminated)
		.reset_req_in5  (1'b0),                            // (terminated)
		.reset_in6      (1'b0),                            // (terminated)
		.reset_req_in6  (1'b0),                            // (terminated)
		.reset_in7      (1'b0),                            // (terminated)
		.reset_req_in7  (1'b0),                            // (terminated)
		.reset_in8      (1'b0),                            // (terminated)
		.reset_req_in8  (1'b0),                            // (terminated)
		.reset_in9      (1'b0),                            // (terminated)
		.reset_req_in9  (1'b0),                            // (terminated)
		.reset_in10     (1'b0),                            // (terminated)
		.reset_req_in10 (1'b0),                            // (terminated)
		.reset_in11     (1'b0),                            // (terminated)
		.reset_req_in11 (1'b0),                            // (terminated)
		.reset_in12     (1'b0),                            // (terminated)
		.reset_req_in12 (1'b0),                            // (terminated)
		.reset_in13     (1'b0),                            // (terminated)
		.reset_req_in13 (1'b0),                            // (terminated)
		.reset_in14     (1'b0),                            // (terminated)
		.reset_req_in14 (1'b0),                            // (terminated)
		.reset_in15     (1'b0),                            // (terminated)
		.reset_req_in15 (1'b0)                             // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),        // reset_in1.reset
		.clk            (altpll_0_c1_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
